package riscv_32_test_pkg;
`include "riscv-tests/rv32ui-p-addi.mem";
`include "riscv-tests/rv32ui-p-add.mem";
`include "riscv-tests/rv32ui-p-andi.mem";
`include "riscv-tests/rv32ui-p-and.mem";
`include "riscv-tests/rv32ui-p-auipc.mem";
`include "riscv-tests/rv32ui-p-beq.mem";
`include "riscv-tests/rv32ui-p-bge.mem";
`include "riscv-tests/rv32ui-p-bgeu.mem";
`include "riscv-tests/rv32ui-p-blt.mem";
`include "riscv-tests/rv32ui-p-bltu.mem";
`include "riscv-tests/rv32ui-p-bne.mem";
`include "riscv-tests/rv32ui-p-fence_i.mem";
`include "riscv-tests/rv32ui-p-jal.mem";
`include "riscv-tests/rv32ui-p-jalr.mem";
`include "riscv-tests/rv32ui-p-lb.mem";
`include "riscv-tests/rv32ui-p-lbu.mem";
`include "riscv-tests/rv32ui-p-lh.mem";
`include "riscv-tests/rv32ui-p-lhu.mem";
`include "riscv-tests/rv32ui-p-lui.mem";
`include "riscv-tests/rv32ui-p-lw.mem";
`include "riscv-tests/rv32ui-p-ori.mem";
`include "riscv-tests/rv32ui-p-or.mem";
`include "riscv-tests/rv32ui-p-sb.mem";
`include "riscv-tests/rv32ui-p-sh.mem";
`include "riscv-tests/rv32ui-p-simple.mem";
`include "riscv-tests/rv32ui-p-slli.mem";
`include "riscv-tests/rv32ui-p-sll.mem";
`include "riscv-tests/rv32ui-p-slti.mem";
`include "riscv-tests/rv32ui-p-sltiu.mem";
`include "riscv-tests/rv32ui-p-slt.mem";
`include "riscv-tests/rv32ui-p-sltu.mem";
`include "riscv-tests/rv32ui-p-srai.mem";
`include "riscv-tests/rv32ui-p-sra.mem";
`include "riscv-tests/rv32ui-p-srli.mem";
`include "riscv-tests/rv32ui-p-srl.mem";
`include "riscv-tests/rv32ui-p-sub.mem";
`include "riscv-tests/rv32ui-p-sw.mem";
`include "riscv-tests/rv32ui-p-xori.mem";
`include "riscv-tests/rv32ui-p-xor.mem";
endpackage
