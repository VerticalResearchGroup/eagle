module l2_cache (
input clk,
input rst_n,
routertollc_request.receiver l2_req,
llctorouter_response.sender  l2_rsp
);


endmodule
