// Tile Operations
`define OP_NOP       0
`define OP_DISPATCH  1
`define OP_COMPLETED 2
